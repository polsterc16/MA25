--
-- VHDL Architecture proj_master_2025_lib.c_006_logic_gate.rtl_xor
--
-- Created:
--          by - Admin.UNKNOWN (LAPTOP-7KFJT032)
--          at - 11:42:58 20.03.2025
--
-- using Mentor Graphics HDL Designer(TM) 2017.1a (Build 5)
--
architecture rtl_xor of c_006_logic_gate is
begin
  out1 <= in1 xor in2;
end architecture rtl_xor;

