--
-- VHDL Architecture proj_master_2025_lib.c_001_binary_counter.rtl
--
-- Created:
--          by - Admin.UNKNOWN (LAPTOP-7KFJT032)
--          at - 08:57:36 11.03.2025
--
-- using Mentor Graphics HDL Designer(TM) 2017.1a (Build 5)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity c_001_binary_counter is
end entity c_001_binary_counter;

--
architecture rtl of c_001_binary_counter is
begin
end architecture rtl;

